module rtl;


endmodule